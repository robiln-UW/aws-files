`ifndef CL_LED_DIP
`define CL_LED_DIP

`define CL_NAME cl_led_dip

`define FPGA_LESS_RST

`endif
